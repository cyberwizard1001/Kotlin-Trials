module orgate(a,b,y);
input a,b;
assign y = a | b;
endmodule
