module and_using_nand(x, y, z);
input a,b;
output c;

nandgate test_gate(c,a,b);


endmodule
