module alu();
